`define C_PCIE_IRQ_CNT  16
`define C_PRJ_SHASUM    0x86b83613
`define C_PRJ_TIMESTAMP 1695192362
`define C_PRJ_VERSION   0x02010001
`define C_TIMESTAMP     1695192362
`define C_VERSION       0x0000002a
