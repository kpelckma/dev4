`define C_DAQ1_CHANNELS_IN_TAB 8
`define C_DAQ2_CHANNELS_IN_TAB 8
`define C_DAQ0_BUF1_OFFSET     1048576
`define C_TRG_CNT              3
`define C_DAQ1_MAX_TRIGGERS    510
`define C_DAQ1_BUF1_OFFSET     5242880
`define C_DAQ2_BUF1_OFFSET     3145728
`define C_DAQ0_TAB_COUNT       1
`define C_DAQ_REGIONS          1
`define C_RTM_TYPE             1
`define C_TIMESTAMP            1695192362
`define C_DAQ1_TAB_COUNT       1
`define C_DAQ2_TAB_COUNT       1
`define C_CHANNEL_WIDTH_BYTES  4
`define C_VERSION              0x02000201
`define C_DAQ0_IS_CONTINUOUS   0
`define C_DAQ0_MAX_SAMPLES     16384
`define C_PRJ_TIMESTAMP        1695192362
`define C_DAQ0_BUF0_OFFSET     0
`define C_DAQ1_IS_CONTINUOUS   0
`define C_DAQ1_MAX_SAMPLES     16384
`define C_DAQ1_BUF0_OFFSET     4194304
`define C_DAQ2_MAX_SAMPLES     16384
`define C_DAQ2_IS_CONTINUOUS   0
`define C_DAQ0_MAX_TRIGGERS    510
`define C_PRJ_VERSION          0x02010001
`define C_DAQ2_BUF0_OFFSET     2097152
`define C_DAQ2_MAX_TRIGGERS    510
`define C_OUT_TRG              3
`define C_PRJ_SHASUM           0x86b83613
`define C_ID                   0x00000002
`define C_DAQ0_CHANNELS_IN_TAB 8
`define C_EXT_TRG              8
