-------------------------------------------------------------------------------
--          ____  _____________  __                                          --
--         / __ \/ ____/ ___/\ \/ /                 _   _   _                --
--        / / / / __/  \__ \  \  /                 / \ / \ / \               --
--       / /_/ / /___ ___/ /  / /               = ( M | S | K )=             --
--      /_____/_____//____/  /_/                   \_/ \_/ \_/               --
--                                                                           --
-------------------------------------------------------------------------------
--! @copyright Copyright 2021 DESY
--! SPDX-License-Identifier: CERN-OHL-W-2.0
-------------------------------------------------------------------------------
--! @date 2022-04-20
--! @author Radoslaw Rybaniec
-------------------------------------------------------------------------------
--! @brief
--! First In First Out buffer, functions package
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package memory_ram is

  
end package memory_ram;
