------------------------------------------------------------------------------
--          ____  _____________  __                                         --
--         / __ \/ ____/ ___/\ \/ /                 _   _   _               --
--        / / / / __/  \__ \  \  /                 / \ / \ / \              --
--       / /_/ / /___ ___/ /  / /               = ( M | S | K )=            --
--      /_____/_____//____/  /_/                   \_/ \_/ \_/              --
--                                                                          --
------------------------------------------------------------------------------
--! @copyright Copyright 2022 DESY
--! SPDX-License-Identifier: CERN-OHL-W-2.0
------------------------------------------------------------------------------
--! @date 2022-04-01
--! @author Lukasz Butkowski  <lukasz.butkowski@desy.de>
------------------------------------------------------------------------------
--! @brief
--! Package with DESY library math components
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package dsp_filter is


end package dsp_filter;
