------------------------------------------------------------------------------
--          ____  _____________  __                                         --
--         / __ \/ ____/ ___/\ \/ /                 _   _   _               --
--        / / / / __/  \__ \  \  /                 / \ / \ / \              --
--       / /_/ / /___ ___/ /  / /               = ( M | S | K )=            --
--      /_____/_____//____/  /_/                   \_/ \_/ \_/              --
--                                                                          --
------------------------------------------------------------------------------
-- @copyright Copyright 2018-2022 DESY
-- SPDX-License-Identifier: CERN-OHL-W-2.0
------------------------------------------------------------------------------
-- @date 2018-10-25/2022-04-04
-- @author Radoslaw Rybaniec
-- @author Lukasz Butkowski <lukasz.butkowski@desy.de>
-- @author Cagil Gumus <cagil.guemues@desy.de>
------------------------------------------------------------------------------
-- @brief
-- i2c sub system for dwc8vm1 rtm module
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;

use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

library desy;
use desy.common_types.all;

library desyrdl;
use desyrdl.pkg_rtm.all;

entity rtm_dwc8vm1_top is
  generic (
    G_CLK_FREQ : natural := 100_000_000);
  port (
    pi_clock : in std_logic;
    pi_reset : in std_logic;

    -- register interface
    pi_s_reg_reset : in  std_logic;
    pi_s_reg : in  t_rtm_m2s;
    po_s_reg : out t_rtm_s2m;
    
    pi_interlock     : in std_logic;   -- interlock generated by application
    po_ext_interlock : out std_logic;  -- external interlock coming into rtm
    -- Zone 3 Signals
    pio_rtm_io_p : inout std_logic_vector(11 downto 0);
    pio_rtm_io_n : inout std_logic_vector(11 downto 0)
  );
end rtm_dwc8vm1_top;

architecture rtl of rtm_dwc8vm1_top is

  signal addrmap_i : t_addrmap_rtm_in;
  signal addrmap_o : t_addrmap_rtm_out;

  signal sig_sdi  : std_logic ;
  signal sig_sdo  : std_logic ;
  signal sig_sdt  : std_logic ;
  signal sig_sci  : std_logic ;
  signal sig_sco  : std_logic ;
  signal sig_sct  : std_logic ;

  signal sig_ext_interlock      : std_logic_vector(0 downto 0); -- external interlock from rtm
  signal sig_ext_interlock_buf  : std_logic_vector(0 downto 0); -- synched external interlock signal from rtm
  signal sig_asych_interlock    : std_logic;
  signal sig_interlock          : std_logic;

  attribute async_reg : string;
  -- designates sig_asych_interlock as receiving asynchronous data
  attribute async_reg of sig_asych_interlock:   signal is "true";
  attribute async_reg of sig_ext_interlock_buf: signal is "true";

begin

  -- ==========================================================================
  ins_desyrdl : entity desyrdl.rtm
  port map (
    pi_clock     => pi_clock,
    pi_reset     => pi_s_reg_reset,
    pi_s_top     => pi_s_reg,
    po_s_top     => po_s_reg,
    pi_addrmap   => addrmap_i,
    po_addrmap   => addrmap_o
  );

  -- ==============================================================================
  blk_rtm_io : block
  begin

    ins_hrl_ibuf_p : iobuf port map (io => pio_rtm_io_p(3), i => sig_sdo, o => sig_sdi, t => "not"(sig_sdt));
    ins_hrl_ibuf_n : iobuf port map (io => pio_rtm_io_n(3), i => sig_sco, o => sig_sci, t => "not"(sig_sct));

    pio_rtm_io_p(10) <= sig_interlock;
    pio_rtm_io_n(10) <= 'Z' ;-- switching to single ended because default application pin constrains are differential
                             -- however on struck this pin is single ended

    inst_ibufds : ibufds
    generic map (
      diff_term => true) -- differential termination
    port map (
      o  => sig_ext_interlock(0),
      i  => pio_rtm_io_p(4),
      ib => pio_rtm_io_n(4)
    );

    po_ext_interlock <= sig_ext_interlock_buf(0);

  end block blk_rtm_io;

  --============================================================================
  -- main RTM logic
  blk_rtm_logic : block
    signal l_adc_a_str  : std_logic;
    signal l_adc_b_str  : std_logic;
    signal l_adc_c_str  : std_logic;
    signal l_adc_d_str  : std_logic;
    signal l_hyt271_trg : std_logic := '0'; -- trigger conversion
    signal timer        : natural := 0;

  begin

    sig_interlock <= addrmap_o.RF_PERMIT.data.data(0) and not pi_interlock;
    addrmap_i.EXT_INTERLOCK.data.data <= sig_ext_interlock;

    -- synching external interlock to improve metastability
    prs_synch_interlock: process(pi_clock, pi_reset)
    begin
      if pi_reset = '1' then
        sig_asych_interlock   <= '0';
        sig_ext_interlock_buf(0) <= '0';
      elsif rising_edge(pi_clock) then
        sig_asych_interlock <= sig_ext_interlock(0);
        sig_ext_interlock_buf(0) <= sig_asych_interlock;
      end if;
    end process;

    -- Periodical readout of the ADC and HYT271 if enabled by the user
    proc_trg:
    process(pi_clock)
    begin
      if rising_edge(pi_clock) then
        if timer >= G_CLK_FREQ then
          l_adc_a_str  <= addrmap_o.ADC_READ_ENA.data.data(0);
          l_adc_b_str  <= addrmap_o.ADC_READ_ENA.data.data(1);
          l_adc_c_str  <= addrmap_o.ADC_READ_ENA.data.data(2);
          l_adc_d_str  <= addrmap_o.ADC_READ_ENA.data.data(3);
          l_hyt271_trg <= addrmap_o.HYT271_READ_ENA.data.data(0);
          timer        <= 0;
        else
          l_adc_a_str  <= '0';
          l_adc_b_str  <= '0';
          l_adc_c_str  <= '0';
          l_adc_d_str  <= '0';
          l_hyt271_trg <= '0';
          timer <= timer + 1;
        end if;
      end if;
    end process;

    ins_i2c_subsys : entity work.i2c_subsys
      generic map (
        G_I2C_CLK_DIV => G_CLK_FREQ/100_000)
      port map (
        pi_reset       => pi_reset,
        pi_clock       => pi_clock,
        po_slow_clk    => open,

        pi_att_val    => addrmap_o.ATT_VAL.data.data,
        pi_att_sel    => addrmap_o.ATT_SEL.data.data,
        pi_att_start  => addrmap_o.ATT_VAL.data.swmod,
        po_att_status => addrmap_i.ATT_STATUS.data.data(0),

        pi_dacab_data => addrmap_o.DACAB.data.data,
        pi_dacab_str  => addrmap_o.DACAB.data.swmod,

        pi_daca_data => addrmap_o.DAC(0).data.data,
        pi_daca_str  => addrmap_o.DAC(0).data.swmod,
        pi_dacb_data => addrmap_o.DAC(1).data.data,
        pi_dacb_str  => addrmap_o.DAC(1).data.swmod,

        po_dac_strobed => open,
        po_dac_status  => addrmap_i.DAC_STATUS.data.data,

        po_adc_a_data => addrmap_i.ADC_A.data.data,
        pi_adc_a_str  => l_adc_a_str,
        po_adc_b_data => addrmap_i.ADC_B.data.data,
        pi_adc_b_str  => l_adc_b_str,
        po_adc_c_data => addrmap_i.ADC_C.data.data,
        pi_adc_c_str  => l_adc_c_str,
        po_adc_d_data => addrmap_i.ADC_D.data.data,
        pi_adc_d_str  => l_adc_d_str,
        po_adc_status => addrmap_i.ADC_STATUS.data.data,

        pi_hyt271_trg  => l_hyt271_trg,
        po_hyt271_humi => addrmap_i.HYT271_HUMI.data.data,
        po_hyt271_temp => addrmap_i.HYT271_TEMP.data.data,
        po_hyt271_done => open,

        pi_sdi => sig_sdi,
        po_sdo => sig_sdo,
        po_sdt => sig_sdt,
        pi_sci => sig_sci,
        po_sco => sig_sco,
        po_sct => sig_sct
      );

  end block blk_rtm_logic;

end rtl;
