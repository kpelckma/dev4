------------------------------------------------------------------------------
--          ____  _____________  __                                         --
--         / __ \/ ____/ ___/\ \/ /                 _   _   _               --
--        / / / / __/  \__ \  \  /                 / \ / \ / \              --
--       / /_/ / /___ ___/ /  / /               = ( M | S | K )=            --
--      /_____/_____//____/  /_/                   \_/ \_/ \_/              --
--                                                                          --
------------------------------------------------------------------------------
--! @copyright Copyright 2023 DESY
--! SPDX-License-Identifier: CERN-OHL-W-2.0
------------------------------------------------------------------------------
--! @date 2023-02-13
--! @author Katharina Schulz  <katharina.schulz@desy.de>
------------------------------------------------------------------------------
--! @brief
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package pkg_config is
  
  constant C_AXI4L_ADDR_WIDTH             : natural := 32;
  constant C_AXI4L_DATA_WIDTH             : natural := 32;

end pkg_config;